// Empty file for now